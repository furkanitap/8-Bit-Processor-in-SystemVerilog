`timescale 1ns / 1ps

module Extend(
    input [5:0] in,
    output [7:0] out
    );
assign out = in; 

endmodule
